`include "mux21_barrel_shifter"
`include "mux41_barrel_shifter"
module barrel_shifter(
	input [7:0]din,
	input [2:0]shamt,
	input LR,
	input AL,
	output [7:0]dout
	);

	
wire w0;
wire w1,w2,w3,w4,w5,w6,w7,w8;
wire w9,w10,w11,w12,w13,w14,w15,w16;
mux21 mux21(.X0(0),.X1(din[7]),.Y(AL),.F(w0));


mux41 m1_31(.X0(din[31]),.X1(w0),.X2(din[31]),.X3(din[30]),.Y({LR,shamt[0]}),.F(w1_31));
mux41 m1_30(.X0(din[30]),.X1(din[31]),.X2(din[30]),.X3(din[29]),.Y({LR,shamt[0]}),.F(w1_30));
mux41 m1_29(.X0(din[29]),.X1(din[30]),.X2(din[29]),.X3(din[28]),.Y({LR,shamt[0]}),.F(w1_29));
mux41 m1_28(.X0(din[28]),.X1(din[29]),.X2(din[28]),.X3(din[27]),.Y({LR,shamt[0]}),.F(w1_28));
mux41 m1_27(.X0(din[27]),.X1(din[28]),.X2(din[27]),.X3(din[26]),.Y({LR,shamt[0]}),.F(w1_27));
mux41 m1_26(.X0(din[26]),.X1(din[27]),.X2(din[26]),.X3(din[25]),.Y({LR,shamt[0]}),.F(w1_26));
mux41 m1_25(.X0(din[25]),.X1(din[26]),.X2(din[25]),.X3(din[24]),.Y({LR,shamt[0]}),.F(w1_25));
mux41 m1_24(.X0(din[24]),.X1(din[25]),.X2(din[24]),.X3(din[23]),.Y({LR,shamt[0]}),.F(w1_24));
mux41 m1_23(.X0(din[23]),.X1(din[24]),.X2(din[23]),.X3(din[22]),.Y({LR,shamt[0]}),.F(w1_23));
mux41 m1_22(.X0(din[22]),.X1(din[23]),.X2(din[22]),.X3(din[21]),.Y({LR,shamt[0]}),.F(w1_22));
mux41 m1_21(.X0(din[21]),.X1(din[22]),.X2(din[21]),.X3(din[20]),.Y({LR,shamt[0]}),.F(w1_21));
mux41 m1_20(.X0(din[20]),.X1(din[21]),.X2(din[20]),.X3(din[19]),.Y({LR,shamt[0]}),.F(w1_20));
mux41 m1_19(.X0(din[19]),.X1(din[20]),.X2(din[19]),.X3(din[18]),.Y({LR,shamt[0]}),.F(w1_19));
mux41 m1_18(.X0(din[18]),.X1(din[19]),.X2(din[18]),.X3(din[17]),.Y({LR,shamt[0]}),.F(w1_18));
mux41 m1_17(.X0(din[17]),.X1(din[18]),.X2(din[17]),.X3(din[16]),.Y({LR,shamt[0]}),.F(w1_17));
mux41 m1_16(.X0(din[16]),.X1(din[17]),.X2(din[16]),.X3(din[15]),.Y({LR,shamt[0]}),.F(w1_16));
mux41 m1_15(.X0(din[15]),.X1(din[16]),.X2(din[15]),.X3(din[14]),.Y({LR,shamt[0]}),.F(w1_15));
mux41 m1_14(.X0(din[14]),.X1(din[15]),.X2(din[14]),.X3(din[13]),.Y({LR,shamt[0]}),.F(w1_14));
mux41 m1_13(.X0(din[13]),.X1(din[14]),.X2(din[13]),.X3(din[12]),.Y({LR,shamt[0]}),.F(w1_13));
mux41 m1_12(.X0(din[12]),.X1(din[13]),.X2(din[12]),.X3(din[11]),.Y({LR,shamt[0]}),.F(w1_12));
mux41 m1_11(.X0(din[11]),.X1(din[12]),.X2(din[11]),.X3(din[10]),.Y({LR,shamt[0]}),.F(w1_11));
mux41 m1_10(.X0(din[10]),.X1(din[11]),.X2(din[10]),.X3(din[9]),.Y({LR,shamt[0]}),.F(w1_10));
mux41 m1_9(.X0(din[9]),.X1(din[10]),.X2(din[9]),.X3(din[8]),.Y({LR,shamt[0]}),.F(w1_9));
mux41 m1_8(.X0(din[8]),.X1(din[9]),.X2(din[8]),.X3(din[7]),.Y({LR,shamt[0]}),.F(w1_8));
mux41 m1_7(.X0(din[7]),.X1(din[8]),.X2(din[7]),.X3(din[6]),.Y({LR,shamt[0]}),.F(w1_7));
mux41 m1_6(.X0(din[6]),.X1(din[7]),.X2(din[6]),.X3(din[5]),.Y({LR,shamt[0]}),.F(w1_6));
mux41 m1_5(.X0(din[5]),.X1(din[6]),.X2(din[5]),.X3(din[4]),.Y({LR,shamt[0]}),.F(w1_5));
mux41 m1_4(.X0(din[4]),.X1(din[5]),.X2(din[4]),.X3(din[3]),.Y({LR,shamt[0]}),.F(w1_4));
mux41 m1_3(.X0(din[3]),.X1(din[4]),.X2(din[3]),.X3(din[2]),.Y({LR,shamt[0]}),.F(w1_3));
mux41 m1_2(.X0(din[2]),.X1(din[3]),.X2(din[2]),.X3(din[1]),.Y({LR,shamt[0]}),.F(w1_2));
mux41 m1_1(.X0(din[1]),.X1(din[2]),.X2(din[1]),.X3(din[0]),.Y({LR,shamt[0]}),.F(w1_1));
mux41 m1_0(.X0(din[0]),.X1(din[1]),.X2(din[0]),.X3(0),.Y({LR,shamt[0]}),.F(w1_0));


mux41 m2_31(.X0(w1_31),.X1(w0),.X2(w1_31),.X3(w1_29),.Y({LR,shamt[1]}),.F(w2_31));
mux41 m2_30(.X0(w1_30),.X1(w0),.X2(w1_30),.X3(w1_28),.Y({LR,shamt[1]}),.F(w2_30));
mux41 m2_29(.X0(w1_29),.X1(w1_31),.X2(w1_29),.X3(w1_27),.Y({LR,shamt[1]}),.F(w2_29));
mux41 m2_28(.X0(w1_28),.X1(w1_30),.X2(w1_28),.X3(w1_26),.Y({LR,shamt[1]}),.F(w2_28));
mux41 m2_27(.X0(w1_27),.X1(w1_29),.X2(w1_27),.X3(w1_25),.Y({LR,shamt[1]}),.F(w2_27));
mux41 m2_26(.X0(w1_26),.X1(w1_28),.X2(w1_26),.X3(w1_24),.Y({LR,shamt[1]}),.F(w2_26));
mux41 m2_25(.X0(w1_25),.X1(w1_27),.X2(w1_25),.X3(w1_23),.Y({LR,shamt[1]}),.F(w2_25));
mux41 m2_24(.X0(w1_24),.X1(w1_26),.X2(w1_24),.X3(w1_22),.Y({LR,shamt[1]}),.F(w2_24));
mux41 m2_23(.X0(w1_23),.X1(w1_25),.X2(w1_23),.X3(w1_21),.Y({LR,shamt[1]}),.F(w2_23));
mux41 m2_22(.X0(w1_22),.X1(w1_24),.X2(w1_22),.X3(w1_20),.Y({LR,shamt[1]}),.F(w2_22));
mux41 m2_21(.X0(w1_21),.X1(w1_23),.X2(w1_21),.X3(w1_19),.Y({LR,shamt[1]}),.F(w2_21));
mux41 m2_20(.X0(w1_20),.X1(w1_22),.X2(w1_20),.X3(w1_18),.Y({LR,shamt[1]}),.F(w2_20));
mux41 m2_19(.X0(w1_19),.X1(w1_21),.X2(w1_19),.X3(w1_17),.Y({LR,shamt[1]}),.F(w2_19));
mux41 m2_18(.X0(w1_18),.X1(w1_20),.X2(w1_18),.X3(w1_16),.Y({LR,shamt[1]}),.F(w2_18));
mux41 m2_17(.X0(w1_17),.X1(w1_19),.X2(w1_17),.X3(w1_15),.Y({LR,shamt[1]}),.F(w2_17));
mux41 m2_16(.X0(w1_16),.X1(w1_18),.X2(w1_16),.X3(w1_14),.Y({LR,shamt[1]}),.F(w2_16));
mux41 m2_15(.X0(w1_15),.X1(w1_17),.X2(w1_15),.X3(w1_13),.Y({LR,shamt[1]}),.F(w2_15));
mux41 m2_14(.X0(w1_14),.X1(w1_16),.X2(w1_14),.X3(w1_12),.Y({LR,shamt[1]}),.F(w2_14));
mux41 m2_13(.X0(w1_13),.X1(w1_15),.X2(w1_13),.X3(w1_11),.Y({LR,shamt[1]}),.F(w2_13));
mux41 m2_12(.X0(w1_12),.X1(w1_14),.X2(w1_12),.X3(w1_10),.Y({LR,shamt[1]}),.F(w2_12));
mux41 m2_11(.X0(w1_11),.X1(w1_13),.X2(w1_11),.X3(w1_9),.Y({LR,shamt[1]}),.F(w2_11));
mux41 m2_10(.X0(w1_10),.X1(w1_12),.X2(w1_10),.X3(w1_8),.Y({LR,shamt[1]}),.F(w2_10));
mux41 m2_9(.X0(w1_9),.X1(w1_11),.X2(w1_9),.X3(1_7),.Y({LR,shamt[1]}),.F(w2_9));
mux41 m2_8(.X0(w1_8),.X1(w1_10),.X2(w1_8),.X3(1_6),.Y({LR,shamt[1]}),.F(w2_8));
mux41 m2_7(.X0(w1_7),.X1(w1_9),.X2(w1_7),.X3(w1_5),.Y({LR,shamt[1]}),.F(w2_7));
mux41 m2_6(.X0(w1_6),.X1(w1_8),.X2(w1_6),.X3(w1_4),.Y({LR,shamt[1]}),.F(w2_6));
mux41 m2_5(.X0(w1_5),.X1(w1_7),.X2(w1_5),.X3(w1_3),.Y({LR,shamt[1]}),.F(w2_5));
mux41 m2_4(.X0(w1_4),.X1(w1_6),.X2(w1_4),.X3(w1_2),.Y({LR,shamt[1]}),.F(w2_4));
mux41 m2_3(.X0(w1_3),.X1(w1_5),.X2(w1_3),.X3(w1_1),.Y({LR,shamt[1]}),.F(w2_3));
mux41 m2_2(.X0(w1_2),.X1(w1_4),.X2(w1_2),.X3(w1_0),.Y({LR,shamt[1]}),.F(w2_2));
mux41 m2_1(.X0(w1_1),.X1(w1_3),.X2(w1_1),.X3(0),.Y({LR,shamt[1]}),.F(w2_1));
mux41 m2_0(.X0(w1_0),.X1(w1_2),.X2(w1_0),.X3(0),.Y({LR,shamt[1]}),.F(w2_0));


mux41 m3_31(.X0(w2_31),.X1(w0),.X2(w2_31),.X3(w2_27),.Y({LR,shamt[2]}),.F(w3_31));
mux41 m3_30(.X0(w2_30),.X1(w0),.X2(w2_30),.X3(w2_26),.Y({LR,shamt[2]}),.F(w3_30));
mux41 m3_29(.X0(w2_29),.X1(w0),.X2(w2_29),.X3(w2_25),.Y({LR,shamt[2]}),.F(w3_29));
mux41 m3_28(.X0(w2_28),.X1(w0),.X2(w2_28),.X3(w2_24),.Y({LR,shamt[2]}),.F(w3_28));
mux41 m3_27(.X0(w2_27),.X1(w2_31),.X2(w2_27),.X3(w2_23),.Y({LR,shamt[2]}),.F(w3_27));
mux41 m3_26(.X0(w2_26),.X1(w2_30),.X2(w2_26),.X3(w2_22),.Y({LR,shamt[2]}),.F(w3_26));
mux41 m3_25(.X0(w2_25),.X1(w2_29),.X2(w2_25),.X3(w2_21),.Y({LR,shamt[2]}),.F(w3_25));
mux41 m3_24(.X0(w2_24),.X1(w2_28),.X2(w2_24),.X3(w2_20),.Y({LR,shamt[2]}),.F(w3_24));
mux41 m3_23(.X0(w2_23),.X1(w2_27),.X2(w2_23),.X3(w2_19),.Y({LR,shamt[2]}),.F(w3_23));
mux41 m3_22(.X0(w2_22),.X1(w2_26),.X2(w2_22),.X3(w2_18),.Y({LR,shamt[2]}),.F(w3_22));
mux41 m3_21(.X0(w2_21),.X1(w2_25),.X2(w2_21),.X3(w2_17),.Y({LR,shamt[2]}),.F(w3_21));
mux41 m3_20(.X0(w2_20),.X1(w2_24),.X2(w2_20),.X3(w2_16),.Y({LR,shamt[2]}),.F(w3_20));
mux41 m3_19(.X0(w2_19),.X1(w2_23),.X2(w2_19),.X3(w2_15),.Y({LR,shamt[2]}),.F(w3_19));
mux41 m3_18(.X0(w2_18),.X1(w2_22),.X2(w2_18),.X3(w2_14),.Y({LR,shamt[2]}),.F(w3_18));
mux41 m3_17(.X0(w2_17),.X1(w2_21),.X2(w2_17),.X3(w2_13),.Y({LR,shamt[2]}),.F(w3_17));
mux41 m3_16(.X0(w2_16),.X1(w2_20),.X2(w2_16),.X3(w2_12),.Y({LR,shamt[2]}),.F(w3_16));
mux41 m3_15(.X0(w2_15),.X1(w2_19),.X2(w2_15),.X3(w2_11),.Y({LR,shamt[2]}),.F(w3_15));
mux41 m3_14(.X0(w2_14),.X1(w2_18),.X2(w2_14),.X3(w2_10),.Y({LR,shamt[2]}),.F(w3_14));
mux41 m3_13(.X0(w2_13),.X1(w2_17),.X2(w2_13),.X3(w2_9),.Y({LR,shamt[2]}),.F(w3_13));
mux41 m3_12(.X0(w2_12),.X1(w2_16),.X2(w2_12),.X3(w2_8),.Y({LR,shamt[2]}),.F(w3_12));
mux41 m3_11(.X0(w2_11),.X1(w2_15),.X2(w2_11),.X3(w2_7),.Y({LR,shamt[2]}),.F(w3_11));
mux41 m3_10(.X0(w2_10),.X1(w2_14),.X2(w2_10),.X3(w2_6),.Y({LR,shamt[2]}),.F(w3_10));
mux41 m3_9(.X0(w2_9),.X1(w2_13),.X2(w2_9),.X3(w2_5),.Y({LR,shamt[2]}),.F(w3_9));
mux41 m3_8(.X0(w2_8),.X1(w2_12),.X2(w2_8),.X3(w2_4),.Y({LR,shamt[2]}),.F(w3_8));
mux41 m3_7(.X0(w2_7),.X1(w2_11),.X2(w2_7),.X3(w2_3),.Y({LR,shamt[2]}),.F(w3_7));
mux41 m3_6(.X0(w2_6),.X1(w2_10),.X2(w2_6),.X3(w2_2),.Y({LR,shamt[2]}),.F(w3_6));
mux41 m3_5(.X0(w2_5),.X1(w2_9),.X2(w2_5),.X3(w2_1),.Y({LR,shamt[2]}),.F(w3_5));
mux41 m2_4(.X0(w2_4),.X1(w2_8),.X2(w2_4),.X3(w2_0),.Y({LR,shamt[2]}),.F(w3_4));
mux41 m3_3(.X0(w2_3),.X1(w2_7),.X2(w2_3),.X3(0),.Y({LR,shamt[2]}),.F(w3_3));
mux41 m3_2(.X0(w2_2),.X1(w2_6),.X2(w2_2),.X3(0),.Y({LR,shamt[2]}),.F(w3_2));
mux41 m3_1(.X0(w2_1),.X1(w2_5),.X2(w2_1),.X3(0),.Y({LR,shamt[2]}),.F(w3_1));
mux41 m3_0(.X0(w2_0),.X1(w2_4),.X2(w2_0),.X3(0),.Y({LR,shamt[2]}),.F(w3_0));


mux41 m4_31(.X0(w3_31),.X1(w0),.X2(w3_31),.X3(w3_23),.Y({LR,shamt[3]}),.F(w4_31));
mux41 m4_30(.X0(w3_30),.X1(w0),.X2(w3_30),.X3(w3_22),.Y({LR,shamt[3]}),.F(w4_30));
mux41 m4_29(.X0(w3_29),.X1(w0),.X2(w3_29),.X3(w3_21),.Y({LR,shamt[3]}),.F(w4_29));
mux41 m4_28(.X0(w3_28),.X1(w0),.X2(w3_28),.X3(w3_20),.Y({LR,shamt[3]}),.F(w4_28));
mux41 m4_27(.X0(w3_27),.X1(w0),.X2(w3_27),.X3(w3_19),.Y({LR,shamt[3]}),.F(w4_27));
mux41 m4_26(.X0(w3_26),.X1(w0),.X2(w3_26),.X3(w3_18),.Y({LR,shamt[3]}),.F(w4_26));
mux41 m4_25(.X0(w3_25),.X1(w0),.X2(w3_25),.X3(w3_17),.Y({LR,shamt[3]}),.F(w4_25));
mux41 m4_24(.X0(w3_24),.X1(w0),.X2(w3_24),.X3(w3_16),.Y({LR,shamt[3]}),.F(w4_24));
mux41 m4_23(.X0(w3_23),.X1(w2_31),.X2(w3_23),.X3(w3_15),.Y({LR,shamt[3]}),.F(w4_23));
mux41 m4_22(.X0(w3_22),.X1(w2_30),.X2(w3_22),.X3(w3_14),.Y({LR,shamt[3]}),.F(w4_22));
mux41 m4_21(.X0(w3_21),.X1(w3_29),.X2(w3_21),.X3(w3_13),.Y({LR,shamt[3]}),.F(w4_21));
mux41 m4_20(.X0(w3_20),.X1(w3_28),.X2(w3_20),.X3(w3_12),.Y({LR,shamt[3]}),.F(w4_20));
mux41 m4_19(.X0(w3_19),.X1(w3_27),.X2(w3_19),.X3(w3_11),.Y({LR,shamt[3]}),.F(w4_19));
mux41 m4_18(.X0(w3_18),.X1(w3_26),.X2(w3_18),.X3(w3_10),.Y({LR,shamt[3]}),.F(w4_18));
mux41 m4_17(.X0(w3_17),.X1(w3_25),.X2(w3_17),.X3(w3_9),.Y({LR,shamt[2]}),.F(w4_17));
mux41 m4_16(.X0(w3_16),.X1(w3_24),.X2(w3_16),.X3(w3_8),.Y({LR,shamt[2]}),.F(w4_16));
mux41 m4_15(.X0(w3_15),.X1(w3_23),.X2(w3_15),.X3(w3_7),.Y({LR,shamt[2]}),.F(w4_15));
mux41 m4_14(.X0(w3_14),.X1(w3_22),.X2(w3_14),.X3(w3_6),.Y({LR,shamt[2]}),.F(w4_14));
mux41 m4_13(.X0(w3_13),.X1(w3_21),.X2(w3_13),.X3(w3_5),.Y({LR,shamt[2]}),.F(w4_13));
mux41 m4_12(.X0(w3_12),.X1(w3_20),.X2(w3_12),.X3(w3_4),.Y({LR,shamt[2]}),.F(w4_12));
mux41 m4_11(.X0(w3_11),.X1(w3_19),.X2(w3_11),.X3(w3_3),.Y({LR,shamt[2]}),.F(w4_11));
mux41 m4_10(.X0(w3_10),.X1(w3_18),.X2(w3_10),.X3(w3_2),.Y({LR,shamt[2]}),.F(w4_10));
mux41 m4_9(.X0(w3_9),.X1(w3_17),.X2(w3_9),.X3(w3_1),.Y({LR,shamt[2]}),.F(w4_9));
mux41 m4_8(.X0(w3_8),.X1(w3_16),.X2(w3_8),.X3(0),.Y({LR,shamt[2]}),.F(w4_8));
mux41 m4_7(.X0(w3_7),.X1(w3_15),.X2(w3_7),.X3(0),.Y({LR,shamt[2]}),.F(w4_7));
mux41 m4_6(.X0(w3_6),.X1(w3_14),.X2(w3_6),.X3(0),.Y({LR,shamt[2]}),.F(w4_6));
mux41 m4_5(.X0(w3_5),.X1(w3_13),.X2(w3_5),.X3(0),.Y({LR,shamt[2]}),.F(w4_5));
mux41 m4_4(.X0(w3_4),.X1(w3_12),.X2(w3_4),.X3(0),.Y({LR,shamt[2]}),.F(w4_4));
mux41 m4_3(.X0(w3_3),.X1(w3_11),.X2(w3_3),.X3(0),.Y({LR,shamt[2]}),.F(w4_3));
mux41 m4_2(.X0(w3_2),.X1(w3_10),.X2(w3_2),.X3(0),.Y({LR,shamt[2]}),.F(w4_2));
mux41 m4_1(.X0(w3_1),.X1(w3_9),.X2(w3_1),.X3(0),.Y({LR,shamt[2]}),.F(w4_1));
mux41 m4_0(.X0(w3_0),.X1(w3_8),.X2(w3_0),.X3(0),.Y({LR,shamt[2]}),.F(w4_0));

mux41 m5_31(.X0(w4_31),.X1(w0),.X2(w4_31),.X3(w4_15),.Y({LR,shamt[4]}),.F(dout[31]));
mux41 m5_30(.X0(w4_30),.X1(w0),.X2(w4_30),.X3(w4_14),.Y({LR,shamt[4]}),.F(dout[30]));
mux41 m5_29(.X0(w4_29),.X1(w0),.X2(w4_29),.X3(w4_13),.Y({LR,shamt[4]}),.F(dout[29]));
mux41 m5_28(.X0(w4_28),.X1(w0),.X2(w4_28),.X3(w4_12),.Y({LR,shamt[4]}),.F(dout[28]));
mux41 m5_27(.X0(w4_27),.X1(w0),.X2(w4_27),.X3(w4_11),.Y({LR,shamt[4]}),.F(dout[27]));
mux41 m5_26(.X0(w4_26),.X1(w0),.X2(w4_26),.X3(w4_10),.Y({LR,shamt[4]}),.F(dout[26]));
mux41 m5_25(.X0(w4_25),.X1(w0),.X2(w4_25),.X3(w4_9),.Y({LR,shamt[4]}),.F(dout[25]));
mux41 m5_24(.X0(w4_24),.X1(w0),.X2(w4_24),.X3(w4_8),.Y({LR,shamt[4]}),.F(dout[24]));
mux41 m5_23(.X0(w4_23),.X1(w0),.X2(w4_23),.X3(w4_7),.Y({LR,shamt[4]}),.F(dout[23]));
mux41 m5_22(.X0(w4_22),.X1(w0),.X2(w4_22),.X3(w4_6),.Y({LR,shamt[4]}),.F(dout[22]));
mux41 m5_21(.X0(w4_21),.X1(w0),.X2(w4_21),.X3(w4_5),.Y({LR,shamt[4]}),.F(dout[21]));
mux41 m5_20(.X0(w4_20),.X1(w0),.X2(w4_20),.X3(w4_4),.Y({LR,shamt[4]}),.F(dout[20]));
mux41 m5_19(.X0(w4_19),.X1(w0),.X2(w4_19),.X3(w4_3),.Y({LR,shamt[4]}),.F(dout[19]));
mux41 m5_18(.X0(w4_18),.X1(w0),.X2(w4_18),.X3(w4_2),.Y({LR,shamt[4]}),.F(dout[18]));
mux41 m5_17(.X0(w4_17),.X1(w0),.X2(w4_17),.X3(w4_1),.Y({LR,shamt[4]}),.F(dout[17]));
mux41 m5_16(.X0(w4_16),.X1(w0),.X2(w4_16),.X3(w4_0),.Y({LR,shamt[4]}),.F(dout[16]));
mux41 m5_15(.X0(w4_15),.X1(w4_31),.X2(w4_15),.X3(0),.Y({LR,shamt[4]}),.F(dout[15]));
mux41 m5_14(.X0(w4_14),.X1(w4_30),.X2(w4_14),.X3(0),.Y({LR,shamt[4]}),.F(dout[14]));
mux41 m5_13(.X0(w4_13),.X1(w4_29),.X2(w4_13),.X3(0),.Y({LR,shamt[4]}),.F(dout[13]));
mux41 m5_12(.X0(w4_12),.X1(w4_28),.X2(w4_12),.X3(0),.Y({LR,shamt[4]}),.F(dout[12]));
mux41 m5_11(.X0(w4_11),.X1(w4_27),.X2(w4_11),.X3(0),.Y({LR,shamt[4]}),.F(dout[11]));
mux41 m5_10(.X0(w4_10),.X1(w4_26),.X2(w4_10),.X3(0),.Y({LR,shamt[4]}),.F(dout[10]));
mux41 m5_9(.X0(w4_9),.X1(w4_25),.X2(w4_9),.X3(0),.Y({LR,shamt[4]}),.F(dout[9]));
mux41 m5_8(.X0(w4_8),.X1(w4_24),.X2(w4_8),.X3(0),.Y({LR,shamt[4]}),.F(dout[8]));
mux41 m5_7(.X0(w4_7),.X1(w4_23),.X2(w4_7),.X3(0),.Y({LR,shamt[4]}),.F(dout[7]));
mux41 m5_6(.X0(w4_6),.X1(w4_22),.X2(w4_6),.X3(0),.Y({LR,shamt[4]}),.F(dout[6]));
mux41 m5_5(.X0(w4_5),.X1(w4_21),.X2(w4_5),.X3(0),.Y({LR,shamt[4]}),.F(dout[5]));
mux41 m5_4(.X0(w4_4),.X1(w4_20),.X2(w4_4),.X3(0),.Y({LR,shamt[4]}),.F(dout[4]));
mux41 m5_3(.X0(w4_3),.X1(w4_19),.X2(w4_3),.X3(0),.Y({LR,shamt[4]}),.F(dout[3]));
mux41 m5_2(.X0(w4_2),.X1(w4_18),.X2(w4_2),.X3(0),.Y({LR,shamt[4]}),.F(dout[2]));
mux41 m5_1(.X0(w4_1),.X1(w4_17),.X2(w4_1),.X3(0),.Y({LR,shamt[4]}),.F(dout[1]));
mux41 m5_0(.X0(w4_0),.X1(w4_16),.X2(w4_0),.X3(0),.Y({LR,shamt[4]}),.F(dout[0]));
endmodule

